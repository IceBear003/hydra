module find_first_one
(
    input [2047:0] data,
    output reg [10:0] cnt = 11'b0
);

reg update_trigger = 1'b0;

always @(data) begin
    
end

always @(data) begin
    
end

endmodule