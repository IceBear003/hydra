module port_wr_frontend(
    input clk,
    input rst_n,

    /*
     * ????????????????
     */
    input wr_sop,
    input wr_eop,
    input wr_vld,
    input [15:0] wr_data,
    output reg pause,

    /*
     * ?????????????????
     * |- xfer_data_vld - xfer_data???????
     * |- xfer_data - ????????????????????
     * |- end_of_packet - ??????????????????????????
     */
    output ready_to_xfer,
    output reg xfer_data_vld,
    output reg [15:0] xfer_data,
    output reg end_of_packet,

    /*
     * ????????????????
     * |- match_suc - ???????????????????????????????
     * |- match_enable - ?????????????
     * |- new_dest_port, new_length - ??????????????????????(????)
     *                                ????????????SRAM????????????????
     */
    input match_suc,
    output reg match_enable,
    output reg [3:0] new_dest_port,
    output reg [2:0] new_prior,
    output reg [8:0] new_length
);

/*
 * wr_state - ?????????????????????:
 * |- 0 - ??????????????(??????wr_eop?????)
 * |- 1 - ?????????????(wr_sop?????)
 * |- 2 - ?????????????(wr_vld??????????)
 * |- 3 - ????????????(????????????????)
 */
reg [1:0] wr_state;

/*
 * xfer_state - ??????????????????????
 * |- 0 - ?????????????
 * |- 1 - ?????????????????????
 * |- 2 - ???????????????(wr_vld??????????????????????????????????????????????????????)
 */
reg [1:0] xfer_state;

/* ????????
 * |- buffer - ?????????????16??64??FIFO??
 * |- wr_ptr - ???????
 * |- xfer_ptr - ???????????????
 * |- end_ptr - ???????????
 */
reg [15:0] buffer [63:0];
reg [5:0] wr_ptr;
wire [5:0] wr_ptr_pls = wr_ptr + 6'd1;
wire [5:0] wr_ptr_plss = wr_ptr + 6'd2;
reg [5:0] xfer_ptr;
wire [5:0] xfer_ptr_pls = xfer_ptr + 6'd1;
reg [6:0] end_ptr;

reg [8:0] wr_length;

always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        wr_state <= 2'd0;
    end else if(wr_state == 2'd0 && wr_sop) begin
        wr_state <= 2'd1;
    end else if(wr_state == 2'd1 && wr_vld) begin
        wr_state <= 2'd2;
    end else if(wr_state == 2'd2 && wr_length == new_length) begin
        wr_state <= 2'd3;
    end else if(wr_state == 2'd3 && wr_eop) begin
        wr_state <= 2'd0; 
    end
end

always @(posedge clk or negedge rst_n) begin
    if(~rst_n) begin
        wr_ptr <= 0;
    end else if(wr_vld) begin
        buffer[wr_ptr] <= wr_data;
        wr_ptr <= wr_ptr + 1;
        if (wr_state == 2'd1) begin
            /* ?????????????????????????????????????????????? */
            new_dest_port <= wr_data[3:0];
            new_length <= wr_data[15:7];
            new_prior <= wr_data[6:4];
            //$display("new_length = %d",wr_data[15:7]);
        end
    end
end

always @(posedge clk) begin
    if(~rst_n) begin
        end_ptr <= 8'hFF;
    end else if(wr_state == 2'd3) begin
        /* ???????????????wr_ptr???????????????????? */
        end_ptr <= wr_ptr;
    end else if(xfer_state == 2'd1 && xfer_ptr_pls == end_ptr) begin
        end_ptr <= 7'd64;
    end
end

always @(posedge clk) begin
    if(wr_state == 2'd0) begin
        wr_length <= 0;
    end else if (wr_vld) begin
        wr_length <= wr_length + 1;
        ////$display("wr_length = %d",wr_length);
    end
end

always @(posedge clk) begin
    if(~rst_n) begin
        match_enable <= 0;
    end else if(wr_vld && wr_state == 2'd1) begin
        /* ????????? */
        match_enable <= 1;
        //$display("1we");
    end else if(match_suc) begin
        /* ???? */
        match_enable <= 0;
    end
end

/* 
 * ???????????A,B?????????
 * ???B????????????????A???????????????????? 
 * ??????????????match_suc????B??????????match_suc????????????
 */
reg pst_match_suc;

always @(posedge clk) begin
    if(~rst_n) begin
        pst_match_suc <= 0;
    end else if(xfer_state == 3'd0) begin
        pst_match_suc <= 0;
    end else if(match_suc) begin
        pst_match_suc <= 1;
    end
end

always @(posedge clk) begin
    if(~rst_n) begin
        xfer_state <= 2'd0;
    end else if(xfer_state == 2'd0 && (match_suc || pst_match_suc)) begin
        /* ?????????????????? */
        xfer_state <= 2'd1;
    end else if(xfer_state == 2'd1 && xfer_ptr_pls == end_ptr) begin
        /* ??????????????????????? */
        xfer_state <= 2'd0;
        //$display("end_ptr = %d",end_ptr);    
    end else if(xfer_state == 2'd1 && xfer_ptr_pls == wr_ptr) begin
        /* ?????????????????????????????? */
        xfer_state <= 2'd2;
    end else if(xfer_state == 2'd2 && xfer_ptr != wr_ptr) begin
        /* ???????????????????????????? */
        xfer_state <= 2'd1;
    end
    //if(xfer_state == 1)
        //$display("xfer_ptr_pls = %d %d %d %d",xfer_ptr_pls,wr_ptr,end_ptr,xfer_state);
end

assign ready_to_xfer = xfer_state == 2'd0 && (match_suc || pst_match_suc);

always @(posedge clk) begin
    if(~rst_n) begin
        end_of_packet <= 0;
    end else if(xfer_state == 2'd1 && xfer_ptr_pls == end_ptr) begin
        /* ??????????????????????????????????? */
        end_of_packet <= 1;
    end else begin
        end_of_packet <= 0;
    end
end

always @(posedge clk) begin
    if(~rst_n) begin
        xfer_ptr <= 0;
        xfer_data_vld <= 0;
    end else if(xfer_state == 2'd1) begin
        xfer_data <= buffer[xfer_ptr];
        xfer_ptr <= xfer_ptr + 1;
        xfer_data_vld <= 1;
    end else begin
        xfer_data_vld <= 0;
    end
end

/*
 * pause - ????????????????????????????????
 *  I - ?????????????????????????????????????????????????????????
 *  II - ???????????????????SRAM????????????????????????????????????????????????????
 */
 always @(posedge clk) begin
    pause <= (wr_ptr_plss == xfer_ptr) ||
             (wr_ptr_pls == xfer_ptr) ||
             (wr_state == 2'd0 && match_enable && ~match_suc);
end

endmodule