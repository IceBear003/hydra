`include "sram.sv"
`include "ecc_encoder.sv"

module sram_interface
(
    input clk,
    input rst_n,

    input [4:0] time_stamp,
    input [4:0] SRAM_IDX,

    /* 写入 */

    input wr_xfer_data_vld,
    input [15:0] wr_xfer_data,
    input wr_end_of_packet,

    output reg [3:0] wr_packet_dest_port,
    output reg [2:0] wr_packet_prior,
    output reg [15:0] wr_packet_head_addr,
    output reg [15:0] wr_packet_tail_addr,
    output reg wr_packet_join_request,
    output reg [5:0] wr_packet_join_time_stamp,

    input concatenate_enable,
    input [10:0] concatenate_head,
    input [15:0] concatenate_tail,

    /* 读出 */

    input rd_page_down,
    input [10:0] rd_page,

    output reg rd_xfer_data_vld,
    output [15:0] rd_xfer_data,
    output [15:0] rd_next_page,
    output [7:0] rd_ecc_code,

    /* 统计 */

    output reg [10:0] free_space
    
    /* SRAM引出，综合用 */
    // ,(*DONT_TOUCH="YES"*) output wr_en,
    // (*DONT_TOUCH="YES"*) output [13:0] wr_addr,
    // (*DONT_TOUCH="YES"*) output [15:0] din,
    
    // (*DONT_TOUCH="YES"*) output rd_en,
    // (*DONT_TOUCH="YES"*) output [13:0] rd_addr,
    // (*DONT_TOUCH="YES"*) input [15:0] dout
);

/******************************************************************************
 *                                重要存储结构                                 *
 ******************************************************************************/

/* ECC编码存储器 */
(* ram_style = "block" *) reg [7:0] ecc_codes [2047:0];
reg [10:0] ec_wr_addr;
wire [7:0] ec_din;
wire [10:0] ec_rd_addr;
reg [7:0] ec_dout;
always @(posedge clk) begin ecc_codes[ec_wr_addr] <= ec_din; end
always @(posedge clk) begin ec_dout <= ecc_codes[ec_rd_addr]; end

/* ECC加码器 */
reg [15:0] ecc_encoder_buffer [7:0];

always @(posedge clk) begin
    if(wr_xfer_data_vld) begin
        if(wr_batch == 0) begin
            /* 页初时清理缓冲，以免脏数据影响ECC计算 */
            ecc_encoder_buffer[1] <= 16'h0000;
            ecc_encoder_buffer[2] <= 16'h0000;
            ecc_encoder_buffer[3] <= 16'h0000;
            ecc_encoder_buffer[4] <= 16'h0000;
            ecc_encoder_buffer[5] <= 16'h0000;
            ecc_encoder_buffer[6] <= 16'h0000;
            ecc_encoder_buffer[7] <= 16'h0000;
        end
        ecc_encoder_buffer[wr_batch] <= wr_xfer_data;
    end
end

always @(posedge clk) begin
    if(wr_batch == 3'd7 && wr_xfer_data_vld || wr_end_of_packet) begin
        /* 页末时准备将结果写入ECC编码存储器 */
        ec_wr_addr <= wr_page;
    end
end

ecc_encoder ecc_encoder( 
    .data_0(ecc_encoder_buffer[0]),
    .data_1(ecc_encoder_buffer[1]),
    .data_2(ecc_encoder_buffer[2]),
    .data_3(ecc_encoder_buffer[3]),
    .data_4(ecc_encoder_buffer[4]),
    .data_5(ecc_encoder_buffer[5]),
    .data_6(ecc_encoder_buffer[6]),
    .data_7(ecc_encoder_buffer[7]),
    .code(ec_din)
);

/* 生成正在读取的页的校验码 (在page_down信号拉高1周期后可视) */
assign ec_rd_addr = rd_page;
assign rd_ecc_code = ec_dout;

/* 跳转表 */
(* ram_style = "block" *) reg [15:0] jump_table [2047:0];
reg [10:0] jt_wr_addr;
reg [15:0] jt_din;
wire [10:0] jt_rd_addr;
reg [15:0] jt_dout;
always @(posedge clk) begin jump_table[jt_wr_addr] <= jt_din; end
always @(posedge clk) begin jt_dout <= jump_table[jt_rd_addr]; end

/* 跳转表拼接 */
always @(posedge clk) begin
    if(concatenate_enable) begin /* 优先进行不同数据包间跳转表的拼接 */
        jt_wr_addr <= concatenate_head;
        jt_din <= concatenate_tail;
    end else if(wr_xfer_data_vld && wr_page != wr_packet_tail_addr[10:0]) begin /* 正常写入时跳转表连接数据包相邻两页 wr_page -> next_page(np_dout) */
        jt_wr_addr <= wr_page;
        jt_din <= {SRAM_IDX, np_dout};
    end
end

/* 生成正在读取的页的下一页的地址 (在page_down信号拉高1周期后可视) */
assign jt_rd_addr = rd_page;
assign rd_next_page = jt_dout;

/* 空闲队列 FIFO结构的RAM */
(* ram_style = "block" *) reg [10:0] null_pages [2047:0];
reg [10:0] np_wr_addr;
reg [10:0] np_din;
wire [10:0] np_rd_addr;
reg [10:0] np_dout;
always @(posedge clk) begin null_pages[np_wr_addr] <= np_din; end
always @(posedge clk) begin np_dout <= null_pages[np_rd_addr]; end

/*
 * np_head_ptr - 空闲队列的头指针
 * np_tail_ptr - 空闲队列的尾指针
 * np_perfusion - 空闲队列的灌注进度
 */
reg [10:0] np_head_ptr;
reg [10:0] np_tail_ptr;
reg [11:0] np_perfusion;

always @(posedge clk) begin
    if(!rst_n) begin 
        np_head_ptr <= 0;
    end if(wr_batch == 0 && wr_xfer_data_vld) begin /* 在一页刚开始的时候弹出顶页 */
        np_head_ptr <= np_head_ptr + 1;
    end
end

assign np_rd_addr = (wr_state == 2'd0 && wr_xfer_data_vld) 
                    ? np_head_ptr + wr_xfer_data[15:10] /* 在数据包刚开始传输时预测数据包尾页地址 */
                    : np_head_ptr; /* 其他时间查询顶部空页地址 */

always @(posedge clk) begin
    if(!rst_n) begin
        np_perfusion <= 0;  /* 灌注从0开始 */
        np_tail_ptr <= 0;
    end else if(rd_page_down) begin /* 回收读出的页 */
        np_tail_ptr <= np_tail_ptr + 1;
        np_wr_addr <= np_tail_ptr;
        np_din <= rd_page;
    end else if(np_perfusion != 12'd2048) begin /* 灌注到2047结束 */
        np_tail_ptr <= np_tail_ptr + 1;
        np_wr_addr <= np_tail_ptr;
        np_din <= np_perfusion;
        np_perfusion <= np_perfusion + 1;
    end
end

/******************************************************************************
 *                                  写入处理                                   *
 ******************************************************************************/

/*
 * 数据包写入状态
 * |- 0 - 无数据包写入
 * |- 1 - 正在写入数据包的第一页
 * |- 2 - 正在写入数据包的后续页
 */
reg [1:0] wr_state;

always @(posedge clk) begin
    if(!rst_n) begin
        wr_state <= 2'd0;
    end else if(wr_state == 2'd0 && wr_xfer_data_vld) begin
        wr_state <= 2'd1;
    end else if(wr_state == 2'd1 && wr_batch == 3'd7 && wr_xfer_data_vld) begin
        wr_state <= 2'd2;
    end else if(wr_state == 2'd2 && wr_end_of_packet) begin
        wr_state <= 2'd0;
    end
end

/* 正在写入的页 */
reg [10:0] wr_page;
/* 在数据包传输完毕之后的第二个周期重新获取新的wr_page，以规避最后一页数据量过少导致的np_dout还未刷新到新的空闲页的问题 */
reg [1:0] regain_wr_page_tick;

always @(posedge clk) begin
    if(!rst_n) begin
        regain_wr_page_tick <= 2'd0;
    end else if(wr_end_of_packet) begin
        regain_wr_page_tick <= 2'd3;
    end else if(regain_wr_page_tick != 0) begin 
        regain_wr_page_tick <= regain_wr_page_tick - 1;
    end
end

always @(posedge clk) begin
    if(!rst_n) begin
        wr_page <= 0;
    end else if((wr_batch == 3'd7 && wr_xfer_data_vld) || regain_wr_page_tick == 2'd1) begin /* 更新wr_page到新页 */
        wr_page <= np_dout;
    end
end

/* 数据包写入切片下标 */
reg [2:0] wr_batch;

always @(posedge clk) begin
    if(!rst_n) begin
        wr_batch <= 0;
    end else if(wr_end_of_packet) begin
        wr_batch <= 0;
    end else if(wr_xfer_data_vld) begin
        wr_batch <= wr_batch + 1;
    end
end

/* 
 * 在数据包刚写入时生成入队请求基本信息
 * |- wr_packet_dest_port - 数据包目的端口
 * |- wr_packet_prior - 数据包优先级
 * |- wr_packet_head_addr - 数据包头地址
 * |- wr_packet_tail_addr - 数据包尾地址
 */
always @(posedge clk) begin
    if(wr_state == 2'd0 && wr_xfer_data_vld) begin
        wr_packet_dest_port <= wr_xfer_data[3:0];
        wr_packet_prior <= wr_xfer_data[6:4];
        wr_packet_head_addr <= {SRAM_IDX, wr_page};
    end
    if(wr_state == 2'd1 && wr_batch == 3'd1) begin
        wr_packet_tail_addr <= {SRAM_IDX, np_dout};
    end
end

/* 在数据包刚写入时发起入队请求 */
always @(posedge clk) begin
    if(wr_state == 2'd0 && wr_xfer_data_vld) begin
        wr_packet_join_request <= 1;
    end else begin
        wr_packet_join_request <= 0;
    end
end

/* 入队请求时间戳 */
always @(posedge clk) begin
    if(~rst_n) begin 
        wr_packet_join_time_stamp <= 6'd32;
    end if(wr_state == 2'd0 && wr_xfer_data_vld) begin
        wr_packet_join_time_stamp <= {1'b0, time_stamp + 5'd1}; /* +1 是为了与主模块中时间序列新插入的时间戳同步 */
    end else if(time_stamp + 5'd1 == wr_packet_join_time_stamp) begin
        wr_packet_join_time_stamp <= 6'd32; /* 32周期后自动还原，防止重复入队 */
    end
end

/******************************************************************************
 *                                  读出处理                                   *
 ******************************************************************************/

reg [3:0] rd_batch; /* 读出切片下标 */
wire [13:0] sram_rd_addr = {rd_page, rd_page_down ? 3'd0 : rd_batch[2:0]}; /* 翻页时，切片下标应为0，其他时刻则为rd_batch */
always @(posedge clk) begin
    rd_xfer_data_vld <= rd_batch != 4'd8 || rd_page_down;
end

always @(posedge clk) begin
    if(~rst_n) begin
        rd_batch <= 4'd8;
    end if(rd_page_down) begin
        rd_batch <= 1; /* 翻页时，下一刻切片下标应为1 */
    end else if(rd_batch != 4'd8) begin
        rd_batch <= rd_batch + 1;
    end
end

/******************************************************************************
 *                                  统计信息                                   *
 ******************************************************************************/

reg [5:0] packet_length;
always @(posedge clk) begin
    if(wr_state == 2'd0 && wr_xfer_data_vld) begin
        packet_length <= wr_xfer_data[15:10] + 1;
    end
end

always @(posedge clk) begin
    if(~rst_n) begin
        free_space <= 11'd2047;
    end else if(wr_packet_join_request && rd_page_down) begin
        free_space <= free_space - packet_length + 1;
    end else if(wr_packet_join_request) begin
        free_space <= free_space - packet_length;
    end else if(rd_page_down) begin
        free_space <= free_space + 1;
    end
end

wire [13:0] sram_wr_addr = {wr_page, wr_batch};

///* SRAM不引出，调试用
sram sram(
    .clk(clk),
    .rst_n(rst_n),
    .wr_en(wr_xfer_data_vld),
    .wr_addr(sram_wr_addr),
    .din(wr_xfer_data),
    .rd_en(rd_page_down || rd_batch != 4'd8),   //仅在需要读取的时候为1，节省SRAM功耗
    .rd_addr(sram_rd_addr),
    .dout(rd_xfer_data)
); 
//*/

/* SRAM引出，综合用 */
// assign wr_en = wr_xfer_data_vld;
// assign wr_addr = sram_wr_addr;
// assign din = wr_xfer_data;
// assign rd_en = rd_page_down || rd_batch != 4'd8;
// assign rd_addr = sram_rd_addr;
// assign rd_xfer_data = dout;

endmodule