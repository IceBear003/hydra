module port_wr_sram_matcher
#(parameter PORT_IDX = 0) /* ?????????????????(0~15) */
(
    input clk,
    input rst_n,

    /*
     * ?????��???
     * |- match_mode - SRAM??????
     *      |- 0 - ?????????
     *      |- 1 - ?????????
     *      |- 2/3 - ??????????
     * |- match_threshold - ???????????????????????????????�ʦ�???????????
     *      |- ????????? ????0
     *      |- ????????? ????16
     *      |- ?????????? ????31
     */
    input [1:0] match_mode,
    input [4:0] match_threshold,

    /* ????????????? */
    input [3:0] new_dest_port,
    input [8:0] new_length,
    input match_enable,
    output reg match_end,

    /*
     * ???????????? 
     * |- viscous - ?????????????
     * |- matching_next_sram - ??????????????SRAM
     * |- matching_best_sram - ???????????SRAM
     */
    input viscous,
    output reg [4:0] matching_next_sram,
    output reg [4:0] matching_best_sram,

    /* 
     * ???��????SRAM????
     * |- accessible - SRAM??????
     * |- free_space - SRAM??????????
     * |- packet_amount - SRAM???��?????????????????
     */
    input accessible,
    input [10:0] free_space,
    input [8:0] packet_amount
);

/* 
 * ?????
 * |- 0 - ��???
 * |- 1 - ?????(?????match_enable???)
 * |- 2 - ??????(??match_end???????)
 */
reg [1:0] state;

/* 
 * ??????
 * |- matching_find - ??????????????SRAM
 * |- matching_tick - ?????????
 * |- matching_sram - ???????????SRAM(matching_next_sram?????)
 * |- max_amount - ???????SRAM??????????????
 */
reg matching_find;
reg [7:0] matching_tick;
reg [4:0] matching_sram;
reg [8:0] max_amount;

/* ?????????
 * |- old_dest_port - ??????????????????
 * |- old_free_space - ????????SRAM???????
 */
reg [3:0] old_dest_port;
reg [10:0] old_free_space;

always @(posedge clk) begin
    if(~rst_n) begin
        state <= 2'd0;
    end else if(state == 2'd0 && match_enable == 1) begin
        if(new_dest_port == old_dest_port && old_free_space >= new_length && viscous) begin
            /* ????????(?????????????SRAM???????????????????)?????????????????? */
            match_end <= 1;
            state <= 2'd2;
            old_free_space <= old_free_space - new_length;
        end else begin
            match_end <= 0;
            state <= 2'd1;
        end
    end else if(state == 2'd1 && matching_find && matching_tick >= match_threshold) begin
        /* ?????????(??????????��??) */
        match_end <= 1;
        state <= 2'd2;
        old_free_space <= free_space - new_length;
        old_dest_port <= new_dest_port;
    end else if(state == 2'd2) begin
        match_end <= 0;
        state <= 2'd0;
    end
end

always @(posedge clk) begin
    if(state == 2'd1) begin
        matching_tick <= matching_tick + 1;
    end else begin
        matching_tick <= 0;
    end
end

/*
 * ???????????????????????SRAM???
 * ?????????????????????????????free_space?????
 *
 * PORT_IDX?????????????????????????????SRAM???????????????
 */
always @(posedge clk) begin
    if(~rst_n) begin
        case(match_mode)
            1: matching_next_sram <= 5'd16 + PORT_IDX;
            default: matching_next_sram <= {PORT_IDX, 1'b0};
        endcase;
    end else begin
        case(match_mode)
            /* ?????????????????2??SRAM??????????? */
            0: matching_next_sram <= matching_next_sram ^ 5'b00001;
            /* ?????????????????1??SRAM??16?�s????SRAM?????????? */
            1: if(matching_next_sram <= 15) matching_next_sram <= matching_next_sram + 16;
               else if(matching_next_sram == 31) matching_next_sram <= {1'b0, PORT_IDX};
               else matching_next_sram <= matching_next_sram + 1;
            /* ??????????????32?�s????SRAM?????????? */
            default: matching_next_sram <= matching_next_sram + 1;
        endcase
    end
end

always @(posedge clk) begin
    matching_sram <= matching_next_sram;
end

always @(posedge clk) begin
    if(state != 2'd1) begin
        matching_find <= 0;
        max_amount <= 0;
    end else if(accessible) begin                   /* ��????? */
    end else if(free_space < new_length) begin      /* ????? */
    end else if(packet_amount >= max_amount) begin  /* ???????? */
        matching_best_sram <= matching_sram;
        max_amount <= packet_amount;
        matching_find <= 1;
    end
end

endmodule