module sram_interface
(

);

endmodule